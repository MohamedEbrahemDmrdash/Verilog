module SBQM(CLK,RESET,PHOTOCELL,TCOUNT,EMPTY,FULL,PCOUNT,WTIME,PCOUNT_7SEG);
input CLK,RESET;
input [1:0]PHOTOCELL;
input [1:0]TCOUNT;
output EMPTY,FULL;
output [2:0]PCOUNT;
output [4:0]WTIME;
output [6:0]PCOUNT_7SEG;
CU controlundit (PHOTOCELL,CLK,RESET,PCOUNT,EMPTY,FULL,EN,UP_DOWN);
COUNTER count  (UP_DOWN,RESET,CLK,EN,PCOUNT);
rom rom1 ({PCOUNT,TCOUNT},WTIME);
sevenSeg pcount(RESET,{1'b0,PCOUNT},PCOUNT_7SEG);
endmodule 